module BattleShip (
    ports
);
    
endmodule